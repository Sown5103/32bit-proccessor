module processor;

endmodule